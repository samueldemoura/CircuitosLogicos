library IEEE; use IEEE.STD_LOGIC_1164.all;

entity tristate is
	port(a:  in  STD_LOGIC_VECTOR(3 downto 0);
		 en: in  STD_LOGIC;
		 y:  out STD_LOGIC_VECTOR(3 downto 0));
end;

architecture synth of tristate is
begin
	y <= "ZZZZ" when en = '0' else a;
end.